// top_mips_single_cycle.sv
