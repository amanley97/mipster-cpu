// alu.sv
