// regfile.sv
