// cu.sv
