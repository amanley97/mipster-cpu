// DataMem.sv
