// pc_register.sv
