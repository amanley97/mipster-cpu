// InstrMem.sv
