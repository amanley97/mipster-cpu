// mips_single_cycle_tb.sv
